module alu_tb;

	alu a0 (
		
	);

endmodule
